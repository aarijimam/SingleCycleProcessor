module PC(index);
input reg index[3:0];
always @(*)
begin

end